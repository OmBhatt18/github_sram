magic
tech sky130A
timestamp 1729280002
<< nwell >>
rect -441 377 -152 519
<< nmos >>
rect -382 210 -367 252
rect -233 210 -218 252
rect -427 69 -385 84
rect -281 69 -239 84
<< pmos >>
rect -382 397 -367 439
rect -233 397 -218 439
<< ndiff >>
rect -422 240 -382 252
rect -422 222 -415 240
rect -398 222 -382 240
rect -422 210 -382 222
rect -367 240 -329 252
rect -367 222 -352 240
rect -335 222 -329 240
rect -367 210 -329 222
rect -273 244 -233 252
rect -273 221 -268 244
rect -251 221 -233 244
rect -273 210 -233 221
rect -218 245 -182 252
rect -218 222 -204 245
rect -187 222 -182 245
rect -218 210 -182 222
rect -427 116 -385 122
rect -427 99 -417 116
rect -396 99 -385 116
rect -427 84 -385 99
rect -281 117 -239 122
rect -281 100 -271 117
rect -250 100 -239 117
rect -281 84 -239 100
rect -427 52 -385 69
rect -427 35 -418 52
rect -397 35 -385 52
rect -281 55 -239 69
rect -427 28 -385 35
rect -281 38 -272 55
rect -251 38 -239 55
rect -281 29 -239 38
<< pdiff >>
rect -422 432 -382 439
rect -422 404 -414 432
rect -397 404 -382 432
rect -422 397 -382 404
rect -367 433 -328 439
rect -367 405 -353 433
rect -336 405 -328 433
rect -367 397 -328 405
rect -273 430 -233 439
rect -273 405 -265 430
rect -248 405 -233 430
rect -273 397 -233 405
rect -218 431 -182 439
rect -218 406 -204 431
rect -187 406 -182 431
rect -218 397 -182 406
<< ndiffc >>
rect -415 222 -398 240
rect -352 222 -335 240
rect -268 221 -251 244
rect -204 222 -187 245
rect -417 99 -396 116
rect -271 100 -250 117
rect -418 35 -397 52
rect -272 38 -251 55
<< pdiffc >>
rect -414 404 -397 432
rect -353 405 -336 433
rect -265 405 -248 430
rect -204 406 -187 431
<< psubdiff >>
rect -281 174 -256 176
rect -421 155 -379 174
rect -356 155 -317 174
rect -294 155 -233 174
rect -281 152 -256 155
<< nsubdiff >>
rect -422 470 -383 494
rect -359 470 -300 494
rect -276 470 -210 494
<< psubdiffcont >>
rect -379 155 -356 174
rect -317 155 -294 174
<< nsubdiffcont >>
rect -383 470 -359 494
rect -300 470 -276 494
<< poly >>
rect -382 439 -367 454
rect -233 439 -218 454
rect -382 362 -367 397
rect -303 364 -272 373
rect -303 362 -296 364
rect -382 347 -296 362
rect -277 347 -272 364
rect -382 252 -367 347
rect -303 338 -272 347
rect -305 304 -273 312
rect -233 304 -218 397
rect -305 287 -298 304
rect -280 289 -218 304
rect -280 287 -273 289
rect -305 279 -273 287
rect -233 252 -218 289
rect -382 197 -367 210
rect -233 197 -218 210
rect -443 69 -427 84
rect -385 69 -281 84
rect -239 69 -226 84
rect -336 42 -321 69
rect -344 34 -313 42
rect -344 17 -337 34
rect -319 17 -313 34
rect -344 9 -313 17
<< polycont >>
rect -296 347 -277 364
rect -298 287 -280 304
rect -337 17 -319 34
<< locali >>
rect -426 494 -210 499
rect -426 493 -383 494
rect -426 469 -415 493
rect -391 470 -383 493
rect -359 470 -300 494
rect -276 493 -210 494
rect -276 470 -269 493
rect -391 469 -269 470
rect -245 469 -210 493
rect -426 463 -210 469
rect -414 439 -397 463
rect -265 439 -248 463
rect -422 432 -389 439
rect -422 404 -414 432
rect -397 404 -389 432
rect -422 397 -389 404
rect -361 433 -328 439
rect -361 405 -353 433
rect -336 405 -328 433
rect -361 397 -328 405
rect -273 430 -240 439
rect -273 405 -265 430
rect -248 405 -240 430
rect -273 397 -240 405
rect -212 431 -182 439
rect -212 406 -204 431
rect -187 406 -182 431
rect -212 397 -182 406
rect -351 329 -334 397
rect -303 364 -272 373
rect -204 364 -187 397
rect -303 347 -296 364
rect -277 347 -187 364
rect -303 338 -272 347
rect -472 312 -334 329
rect -472 114 -455 312
rect -351 304 -334 312
rect -305 304 -273 312
rect -351 287 -298 304
rect -280 287 -273 304
rect -351 252 -334 287
rect -305 279 -273 287
rect -204 252 -187 347
rect -422 240 -391 252
rect -422 222 -415 240
rect -398 222 -391 240
rect -422 210 -391 222
rect -360 240 -329 252
rect -360 222 -352 240
rect -335 222 -329 240
rect -360 210 -329 222
rect -273 244 -242 252
rect -273 221 -268 244
rect -251 221 -242 244
rect -273 210 -242 221
rect -211 245 -182 252
rect -211 222 -204 245
rect -187 222 -182 245
rect -211 210 -182 222
rect -408 182 -391 210
rect -267 187 -250 210
rect -267 182 -233 187
rect -433 177 -233 182
rect -433 153 -414 177
rect -389 176 -233 177
rect -389 174 -276 176
rect -389 155 -379 174
rect -356 155 -317 174
rect -294 155 -276 174
rect -389 153 -276 155
rect -433 152 -276 153
rect -251 152 -233 176
rect -433 148 -233 152
rect -427 116 -385 122
rect -427 114 -417 116
rect -472 99 -417 114
rect -396 99 -385 116
rect -472 97 -385 99
rect -427 92 -385 97
rect -281 120 -239 122
rect -203 120 -186 210
rect -281 117 -186 120
rect -281 100 -271 117
rect -250 103 -186 117
rect -250 100 -239 103
rect -281 95 -239 100
rect -427 52 -385 58
rect -427 48 -418 52
rect -454 35 -418 48
rect -397 35 -385 52
rect -281 55 -239 61
rect -454 31 -385 35
rect -427 28 -385 31
rect -344 34 -313 42
rect -344 17 -337 34
rect -319 17 -313 34
rect -281 38 -272 55
rect -251 54 -239 55
rect -251 38 -207 54
rect -281 37 -207 38
rect -281 29 -239 37
rect -344 9 -313 17
rect -337 -13 -319 9
<< viali >>
rect -415 469 -391 493
rect -269 469 -245 493
rect -414 153 -389 177
rect -276 152 -251 176
<< metal1 >>
rect -432 493 -210 506
rect -432 469 -415 493
rect -391 469 -269 493
rect -245 469 -210 493
rect -432 459 -210 469
rect -433 177 -233 187
rect -433 153 -414 177
rect -389 176 -233 177
rect -389 153 -276 176
rect -433 152 -276 153
rect -251 152 -233 176
rect -433 145 -233 152
<< labels >>
flabel metal1 -355 465 -301 494 0 FreeSans 152 0 0 0 vdd
flabel locali -216 349 -187 363 0 FreeSans 104 0 0 0 qbar
flabel locali -449 313 -425 328 0 FreeSans 104 0 0 0 q
flabel metal1 -354 157 -319 174 0 FreeSans 120 0 0 0 gnd
flabel locali -336 -7 -321 7 0 FreeSans 72 0 0 0 wl
flabel locali -232 37 -216 54 0 FreeSans 40 0 0 0 blbar_noconn
flabel locali -453 31 -440 48 0 FreeSans 40 0 0 0 bl_noconn
<< end >>
