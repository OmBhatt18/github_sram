magic
tech sky130A
timestamp 1729278784
<< end >>
