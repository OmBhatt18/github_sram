magic
tech sky130A
timestamp 1729279007
<< nwell >>
rect -30 198 127 418
rect 255 176 535 430
rect 255 175 457 176
<< nmos >>
rect 59 537 74 579
rect 320 537 335 579
rect 464 537 479 579
rect 605 537 620 579
rect 59 41 74 83
rect 312 40 327 82
rect 464 40 479 82
rect 603 40 618 82
<< pmos >>
rect 59 358 74 400
rect 59 216 74 258
rect 320 368 335 410
rect 464 368 479 410
rect 312 195 327 237
rect 464 195 479 237
<< ndiff >>
rect 20 570 59 579
rect 20 553 26 570
rect 43 553 59 570
rect 20 537 59 553
rect 74 568 114 579
rect 74 551 88 568
rect 105 551 114 568
rect 74 537 114 551
rect 280 568 320 579
rect 280 549 284 568
rect 303 549 320 568
rect 280 537 320 549
rect 335 568 376 579
rect 335 549 351 568
rect 370 549 376 568
rect 335 537 376 549
rect 417 566 464 579
rect 417 547 423 566
rect 442 547 464 566
rect 417 537 464 547
rect 479 569 535 579
rect 479 550 509 569
rect 528 550 535 569
rect 479 537 535 550
rect 564 567 605 579
rect 564 548 569 567
rect 588 548 605 567
rect 564 537 605 548
rect 620 565 661 579
rect 620 546 636 565
rect 655 546 661 565
rect 620 537 661 546
rect 20 67 59 83
rect 20 50 26 67
rect 43 50 59 67
rect 20 41 59 50
rect 74 69 114 83
rect 74 52 88 69
rect 105 52 114 69
rect 74 41 114 52
rect 274 73 312 82
rect 274 51 279 73
rect 297 51 312 73
rect 274 40 312 51
rect 327 72 365 82
rect 327 50 343 72
rect 361 50 365 72
rect 327 40 365 50
rect 420 72 464 82
rect 420 50 426 72
rect 444 50 464 72
rect 420 40 464 50
rect 479 73 523 82
rect 479 51 495 73
rect 513 51 523 73
rect 479 40 523 51
rect 561 71 603 82
rect 561 51 567 71
rect 584 51 603 71
rect 561 40 603 51
rect 618 74 663 82
rect 618 52 641 74
rect 659 52 663 74
rect 618 40 663 52
<< pdiff >>
rect 24 391 59 400
rect 24 368 29 391
rect 46 368 59 391
rect 24 358 59 368
rect 74 391 109 400
rect 74 368 88 391
rect 105 368 109 391
rect 74 358 109 368
rect 24 248 59 258
rect 24 225 29 248
rect 46 225 59 248
rect 24 216 59 225
rect 74 248 109 258
rect 74 225 88 248
rect 105 225 109 248
rect 74 216 109 225
rect 285 402 320 410
rect 285 379 289 402
rect 306 379 320 402
rect 285 368 320 379
rect 335 399 370 410
rect 335 376 348 399
rect 365 376 370 399
rect 335 368 370 376
rect 427 402 464 410
rect 427 379 434 402
rect 451 379 464 402
rect 427 368 464 379
rect 479 402 516 410
rect 479 379 494 402
rect 511 379 516 402
rect 479 368 516 379
rect 279 226 312 237
rect 279 203 283 226
rect 300 203 312 226
rect 279 195 312 203
rect 327 229 360 237
rect 327 206 336 229
rect 353 206 360 229
rect 327 195 360 206
rect 427 226 464 237
rect 427 203 433 226
rect 450 203 464 226
rect 427 195 464 203
rect 479 226 516 237
rect 479 203 494 226
rect 511 203 516 226
rect 479 195 516 203
<< ndiffc >>
rect 26 553 43 570
rect 88 551 105 568
rect 284 549 303 568
rect 351 549 370 568
rect 423 547 442 566
rect 509 550 528 569
rect 569 548 588 567
rect 636 546 655 565
rect 26 50 43 67
rect 88 52 105 69
rect 279 51 297 73
rect 343 50 361 72
rect 426 50 444 72
rect 495 51 513 73
rect 567 51 584 71
rect 641 52 659 74
<< pdiffc >>
rect 29 368 46 391
rect 88 368 105 391
rect 29 225 46 248
rect 88 225 105 248
rect 289 379 306 402
rect 348 376 365 399
rect 434 379 451 402
rect 494 379 511 402
rect 283 203 300 226
rect 336 206 353 229
rect 433 203 450 226
rect 494 203 511 226
<< psubdiff >>
rect 2 616 56 642
rect 87 616 317 642
rect 348 616 453 642
rect 484 616 553 642
rect 584 616 611 642
rect 266 615 286 616
rect 2 -22 56 4
rect 87 -22 141 4
rect 347 3 413 12
rect 509 3 528 10
rect 257 -23 311 3
rect 342 -23 453 3
rect 484 -23 533 3
rect 564 -23 608 3
rect 347 -24 413 -23
<< nsubdiff >>
rect 22 304 41 305
rect 2 285 45 304
rect 68 285 109 304
rect 273 286 287 305
rect 304 286 331 305
<< psubdiffcont >>
rect 56 616 87 642
rect 317 616 348 642
rect 453 616 484 642
rect 553 616 584 642
rect 56 -22 87 4
rect 311 -23 342 3
rect 453 -23 484 3
rect 533 -23 564 3
<< nsubdiffcont >>
rect 45 285 68 304
rect 287 286 304 305
<< poly >>
rect 59 579 74 592
rect 320 579 335 592
rect 464 579 479 592
rect 605 579 620 592
rect 59 452 74 537
rect 232 506 270 516
rect 320 506 335 537
rect 232 505 335 506
rect 232 486 242 505
rect 260 491 335 505
rect 260 486 270 491
rect 232 478 270 486
rect 59 437 175 452
rect 59 400 74 437
rect 59 345 74 358
rect 59 258 74 271
rect 59 169 74 216
rect -24 159 74 169
rect -24 137 -17 159
rect 3 137 74 159
rect 160 152 175 437
rect 320 410 335 491
rect 464 410 479 537
rect 605 512 620 537
rect 596 504 634 512
rect 596 485 606 504
rect 624 485 634 504
rect 596 474 634 485
rect 320 355 335 368
rect 464 317 479 368
rect 561 320 597 332
rect 561 317 568 320
rect 464 302 568 317
rect 312 237 327 250
rect 464 237 479 302
rect 561 297 568 302
rect 588 297 597 320
rect 561 285 597 297
rect -24 127 74 137
rect 59 83 74 127
rect 152 142 190 152
rect 152 123 160 142
rect 178 139 190 142
rect 312 139 327 195
rect 178 124 327 139
rect 178 123 190 124
rect 152 114 190 123
rect 312 82 327 124
rect 464 82 479 195
rect 587 150 625 158
rect 587 131 597 150
rect 615 131 625 150
rect 587 120 625 131
rect 603 82 618 120
rect 59 28 74 41
rect 312 27 327 40
rect 464 27 479 40
rect 603 27 618 40
<< polycont >>
rect 242 486 260 505
rect -17 137 3 159
rect 606 485 624 504
rect 568 297 588 320
rect 160 123 178 142
rect 597 131 615 150
<< locali >>
rect -5 642 612 643
rect -5 616 56 642
rect 87 635 317 642
rect 87 616 266 635
rect 286 616 317 635
rect 348 616 453 642
rect 484 636 553 642
rect 484 617 517 636
rect 537 617 553 636
rect 484 616 553 617
rect 584 636 612 642
rect 584 617 590 636
rect 610 617 612 636
rect 584 616 612 617
rect -5 614 612 616
rect 27 579 44 614
rect 286 579 304 614
rect 423 579 440 614
rect 569 579 586 614
rect 20 570 52 579
rect 20 553 26 570
rect 43 553 52 570
rect 20 543 52 553
rect 82 568 114 579
rect 82 551 88 568
rect 105 551 114 568
rect 82 543 114 551
rect 280 568 309 579
rect 280 549 284 568
rect 303 549 309 568
rect 89 506 106 543
rect 280 537 309 549
rect 347 568 376 579
rect 347 549 351 568
rect 370 549 376 568
rect 347 537 376 549
rect 417 566 446 579
rect 417 547 423 566
rect 442 547 446 566
rect 417 537 446 547
rect 502 569 531 579
rect 502 550 509 569
rect 528 550 531 569
rect 502 537 531 550
rect 564 567 593 579
rect 564 548 569 567
rect 588 548 593 567
rect 564 537 593 548
rect 632 565 661 579
rect 632 546 636 565
rect 655 563 661 565
rect 655 546 687 563
rect 704 546 707 563
rect 632 537 661 546
rect 232 506 270 516
rect 89 505 270 506
rect 89 489 242 505
rect 89 399 106 489
rect 232 486 242 489
rect 260 486 270 505
rect 232 478 270 486
rect 353 502 370 537
rect 507 502 524 537
rect 596 504 634 512
rect 596 502 606 504
rect 353 485 606 502
rect 624 485 634 504
rect 495 410 512 485
rect 596 474 634 485
rect 285 402 312 410
rect 24 391 51 399
rect 24 368 29 391
rect 46 368 51 391
rect 24 358 51 368
rect 82 391 109 399
rect 82 368 88 391
rect 105 368 109 391
rect 285 379 289 402
rect 306 379 312 402
rect 285 369 312 379
rect 343 399 370 410
rect 343 376 348 399
rect 365 398 370 399
rect 427 402 454 410
rect 427 398 434 402
rect 365 381 434 398
rect 365 376 370 381
rect 82 358 109 368
rect 28 307 45 358
rect 292 308 309 369
rect 343 368 370 376
rect 427 379 434 381
rect 451 379 454 402
rect 427 368 454 379
rect 489 402 516 410
rect 489 379 494 402
rect 511 379 516 402
rect 489 369 516 379
rect 561 320 597 332
rect -3 281 0 307
rect 21 304 91 307
rect 21 285 45 304
rect 68 285 91 304
rect 21 281 91 285
rect 112 281 116 307
rect 273 305 348 308
rect 273 286 287 305
rect 304 302 348 305
rect 304 286 324 302
rect 273 285 324 286
rect 341 285 348 302
rect 561 297 568 320
rect 588 318 597 320
rect 588 301 614 318
rect 588 297 597 301
rect 561 285 597 297
rect 273 282 348 285
rect 28 258 45 281
rect 24 248 51 258
rect 24 225 29 248
rect 46 225 51 248
rect 24 217 51 225
rect 82 248 109 258
rect 82 225 88 248
rect 105 225 109 248
rect 283 236 300 282
rect 82 217 109 225
rect 279 226 306 236
rect -24 159 11 169
rect -24 154 -17 159
rect -45 137 -17 154
rect 3 137 11 159
rect -24 127 11 137
rect 89 141 106 217
rect 279 203 283 226
rect 300 203 306 226
rect 279 195 306 203
rect 333 229 360 237
rect 333 206 336 229
rect 353 226 360 229
rect 427 226 454 237
rect 353 209 433 226
rect 353 206 360 209
rect 333 195 360 206
rect 427 203 433 209
rect 450 203 454 226
rect 427 195 454 203
rect 489 226 516 236
rect 489 203 494 226
rect 511 203 516 226
rect 489 195 516 203
rect 152 142 190 152
rect 495 147 512 195
rect 587 150 625 158
rect 587 147 597 150
rect 152 141 160 142
rect 89 124 160 141
rect 89 77 106 124
rect 152 123 160 124
rect 178 123 190 142
rect 152 114 190 123
rect 343 131 597 147
rect 615 131 625 150
rect 343 130 625 131
rect 343 82 360 130
rect 495 82 512 130
rect 587 120 625 130
rect 20 67 52 77
rect 20 50 26 67
rect 43 50 52 67
rect 20 41 52 50
rect 82 69 114 77
rect 82 52 88 69
rect 105 52 114 69
rect 82 41 114 52
rect 274 73 303 82
rect 274 51 279 73
rect 297 51 303 73
rect 27 12 44 41
rect 274 40 303 51
rect 336 72 365 82
rect 336 50 343 72
rect 361 50 365 72
rect 336 40 365 50
rect 420 72 449 82
rect 420 50 426 72
rect 444 50 449 72
rect 420 40 449 50
rect 489 73 518 82
rect 489 51 495 73
rect 513 51 518 73
rect 489 40 518 51
rect 561 71 592 82
rect 561 51 567 71
rect 584 51 592 71
rect 561 40 592 51
rect 632 74 663 82
rect 632 52 641 74
rect 659 68 663 74
rect 659 52 691 68
rect 632 51 691 52
rect 632 40 663 51
rect -5 11 224 12
rect 280 11 298 40
rect 424 12 441 40
rect 343 11 450 12
rect 496 11 513 12
rect 570 11 587 40
rect -5 4 626 11
rect -5 -13 24 4
rect 41 -13 56 4
rect -5 -22 56 -13
rect 87 3 626 4
rect 87 2 311 3
rect 87 -15 260 2
rect 277 -15 311 2
rect 87 -22 311 -15
rect -5 -23 311 -22
rect 342 0 453 3
rect 342 -17 388 0
rect 405 -17 453 0
rect 342 -23 453 -17
rect 484 -23 533 3
rect 564 -23 577 3
rect 608 -23 626 3
rect 248 -24 626 -23
<< viali >>
rect 266 616 286 635
rect 517 617 537 636
rect 590 617 610 636
rect 687 546 704 563
rect 0 281 21 307
rect 91 281 112 307
rect 324 285 341 302
rect 691 51 708 68
rect 24 -13 41 4
rect 260 -15 277 2
rect 388 -17 405 0
rect 577 -23 608 3
<< metal1 >>
rect -7 636 614 645
rect -7 635 517 636
rect -7 616 266 635
rect 286 617 517 635
rect 537 617 590 636
rect 610 617 614 636
rect 286 616 614 617
rect -7 607 614 616
rect 661 563 710 571
rect 661 546 687 563
rect 704 546 710 563
rect 661 540 710 546
rect -12 307 120 315
rect -12 281 0 307
rect 21 281 91 307
rect 112 281 120 307
rect -12 274 120 281
rect 255 302 348 316
rect 255 285 324 302
rect 341 285 348 302
rect 255 275 348 285
rect 663 68 713 74
rect 663 51 691 68
rect 708 51 713 68
rect 663 46 713 51
rect 699 45 713 46
rect -15 12 44 13
rect -15 4 626 12
rect -15 -13 24 4
rect 41 3 626 4
rect 41 2 577 3
rect 41 -13 260 2
rect -15 -15 260 -13
rect 277 0 577 2
rect 277 -15 388 0
rect -15 -17 388 -15
rect 405 -17 577 0
rect -15 -23 577 -17
rect 608 -23 626 3
rect -15 -32 626 -23
<< labels >>
flabel locali 108 124 131 140 0 FreeSans 80 0 0 0 dinb
flabel metal1 24 283 43 300 0 FreeSans 72 270 0 0 vdd
flabel metal1 307 285 320 302 0 FreeSans 72 270 0 0 vdd
flabel metal1 359 615 413 642 0 FreeSans 152 0 0 0 gnd
flabel metal1 94 -22 141 4 0 FreeSans 152 0 0 0 gnd
flabel locali 91 490 146 505 0 FreeSans 152 0 0 0 dinbb
flabel locali -44 138 -25 153 0 FreeSans 120 0 0 0 din
flabel locali 504 131 545 147 0 FreeSans 144 0 0 0 out1
flabel locali 507 486 539 502 0 FreeSans 144 0 0 0 out2
flabel metal1 663 547 686 563 0 FreeSans 120 0 0 0 bl
flabel metal1 666 53 688 67 0 FreeSans 96 0 0 0 blbar
flabel locali 375 210 405 225 0 FreeSans 120 0 0 0 4
flabel locali 379 382 407 397 0 FreeSans 120 0 0 0 5
flabel locali 599 303 612 315 0 FreeSans 88 0 0 0 wen
<< end >>
