* SPICE3 file created from cell_6t.ext - technology: sky130A
.SUBCKT cell_1rw bl br wl vdd gnd
X0 q qbar gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.168 ps=1.64 w=0.42 l=0.15
X1 q qbar vdd vdd sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.62 as=0.168 ps=1.64 w=0.42 l=0.15
X2 q wl bl gnd sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.1722 ps=1.66 w=0.42 l=0.15
X3 qbar wl br gnd sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.168 ps=1.64 w=0.42 l=0.15
X4 qbar q gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.168 ps=1.64 w=0.42 l=0.15
X5 qbar q vdd vdd sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.62 as=0.168 ps=1.64 w=0.42 l=0.15

.ENDS
