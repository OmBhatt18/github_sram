magic
tech sky130A
timestamp 1729324531
<< nwell >>
rect 559 177 843 319
<< nmos >>
rect 618 10 633 52
rect 767 10 782 52
rect 573 -131 615 -116
rect 719 -131 761 -116
<< pmos >>
rect 618 197 633 239
rect 767 197 782 239
<< ndiff >>
rect 578 40 618 52
rect 578 22 585 40
rect 602 22 618 40
rect 578 10 618 22
rect 633 40 671 52
rect 633 22 648 40
rect 665 22 671 40
rect 633 10 671 22
rect 727 44 767 52
rect 727 21 732 44
rect 749 21 767 44
rect 727 10 767 21
rect 782 45 820 52
rect 782 22 796 45
rect 813 22 820 45
rect 782 10 820 22
rect 573 -84 615 -78
rect 573 -101 583 -84
rect 604 -101 615 -84
rect 573 -116 615 -101
rect 719 -83 761 -78
rect 719 -100 729 -83
rect 750 -100 761 -83
rect 719 -116 761 -100
rect 573 -148 615 -131
rect 573 -165 582 -148
rect 603 -165 615 -148
rect 719 -145 761 -131
rect 573 -172 615 -165
rect 719 -162 728 -145
rect 749 -162 761 -145
rect 719 -171 761 -162
<< pdiff >>
rect 578 232 618 239
rect 578 204 586 232
rect 603 204 618 232
rect 578 197 618 204
rect 633 233 672 239
rect 633 205 647 233
rect 664 205 672 233
rect 633 197 672 205
rect 727 230 767 239
rect 727 205 735 230
rect 752 205 767 230
rect 727 197 767 205
rect 782 231 821 239
rect 782 206 796 231
rect 813 206 821 231
rect 782 197 821 206
<< ndiffc >>
rect 585 22 602 40
rect 648 22 665 40
rect 732 21 749 44
rect 796 22 813 45
rect 583 -101 604 -84
rect 729 -100 750 -83
rect 582 -165 603 -148
rect 728 -162 749 -145
<< pdiffc >>
rect 586 204 603 232
rect 647 205 664 233
rect 735 205 752 230
rect 796 206 813 231
<< psubdiff >>
rect 719 -26 744 -24
rect 579 -45 621 -26
rect 644 -45 683 -26
rect 706 -45 767 -26
rect 719 -48 744 -45
<< nsubdiff >>
rect 578 270 617 294
rect 641 270 700 294
rect 724 270 790 294
<< psubdiffcont >>
rect 621 -45 644 -26
rect 683 -45 706 -26
<< nsubdiffcont >>
rect 617 270 641 294
rect 700 270 724 294
<< poly >>
rect 618 239 633 254
rect 767 239 782 254
rect 618 162 633 197
rect 697 164 728 173
rect 697 162 704 164
rect 618 147 704 162
rect 723 147 728 164
rect 618 52 633 147
rect 697 138 728 147
rect 695 104 727 112
rect 767 104 782 197
rect 695 87 702 104
rect 720 89 782 104
rect 720 87 727 89
rect 695 79 727 87
rect 767 52 782 89
rect 618 -3 633 10
rect 767 -3 782 10
rect 557 -131 573 -116
rect 615 -131 719 -116
rect 761 -131 774 -116
rect 664 -158 679 -131
rect 656 -166 687 -158
rect 656 -183 663 -166
rect 681 -183 687 -166
rect 656 -191 687 -183
<< polycont >>
rect 704 147 723 164
rect 702 87 720 104
rect 663 -183 681 -166
<< locali >>
rect 574 294 790 299
rect 574 293 617 294
rect 574 269 585 293
rect 609 270 617 293
rect 641 270 700 294
rect 724 293 790 294
rect 724 270 731 293
rect 609 269 731 270
rect 755 269 790 293
rect 574 263 790 269
rect 586 239 603 263
rect 735 239 752 263
rect 578 232 611 239
rect 578 204 586 232
rect 603 204 611 232
rect 578 197 611 204
rect 639 233 672 239
rect 639 205 647 233
rect 664 205 672 233
rect 639 197 672 205
rect 727 230 760 239
rect 727 205 735 230
rect 752 205 760 230
rect 727 197 760 205
rect 788 231 821 239
rect 788 206 796 231
rect 813 206 821 231
rect 788 197 821 206
rect 649 129 666 197
rect 697 164 728 173
rect 796 164 813 197
rect 697 147 704 164
rect 723 147 813 164
rect 697 138 728 147
rect 528 112 666 129
rect 528 -86 545 112
rect 649 104 666 112
rect 695 104 727 112
rect 649 87 702 104
rect 720 87 727 104
rect 649 52 666 87
rect 695 79 727 87
rect 796 52 813 147
rect 578 40 609 52
rect 578 22 585 40
rect 602 22 609 40
rect 578 10 609 22
rect 640 40 671 52
rect 640 22 648 40
rect 665 22 671 40
rect 640 10 671 22
rect 727 44 758 52
rect 727 21 732 44
rect 749 21 758 44
rect 727 10 758 21
rect 789 45 820 52
rect 789 22 796 45
rect 813 22 820 45
rect 789 10 820 22
rect 592 -18 609 10
rect 733 -13 750 10
rect 733 -18 767 -13
rect 567 -23 767 -18
rect 567 -47 586 -23
rect 611 -24 767 -23
rect 611 -26 724 -24
rect 611 -45 621 -26
rect 644 -45 683 -26
rect 706 -45 724 -26
rect 611 -47 724 -45
rect 567 -48 724 -47
rect 749 -48 767 -24
rect 567 -52 767 -48
rect 573 -84 615 -78
rect 573 -86 583 -84
rect 528 -101 583 -86
rect 604 -101 615 -84
rect 528 -103 615 -101
rect 573 -108 615 -103
rect 719 -80 761 -78
rect 797 -80 814 10
rect 719 -83 814 -80
rect 719 -100 729 -83
rect 750 -97 814 -83
rect 750 -100 761 -97
rect 719 -105 761 -100
rect 518 -151 543 -142
rect 518 -169 523 -151
rect 540 -152 543 -151
rect 573 -148 615 -142
rect 573 -152 582 -148
rect 540 -165 582 -152
rect 603 -165 615 -148
rect 719 -145 761 -139
rect 540 -169 615 -165
rect 518 -179 543 -169
rect 573 -172 615 -169
rect 656 -166 687 -158
rect 656 -183 663 -166
rect 681 -183 687 -166
rect 719 -162 728 -145
rect 749 -146 761 -145
rect 825 -145 850 -135
rect 825 -146 829 -145
rect 749 -162 829 -146
rect 719 -163 829 -162
rect 846 -163 850 -145
rect 719 -171 761 -163
rect 825 -172 850 -163
rect 656 -191 687 -183
rect 663 -213 681 -191
<< viali >>
rect 585 269 609 293
rect 731 269 755 293
rect 586 -47 611 -23
rect 724 -48 749 -24
rect 523 -169 540 -151
rect 829 -163 846 -145
<< metal1 >>
rect 517 -151 544 331
rect 568 293 790 306
rect 568 269 585 293
rect 609 269 731 293
rect 755 269 790 293
rect 568 259 790 269
rect 567 -23 767 -13
rect 567 -47 586 -23
rect 611 -24 767 -23
rect 611 -47 724 -24
rect 567 -48 724 -47
rect 749 -48 767 -24
rect 567 -55 767 -48
rect 517 -169 523 -151
rect 540 -152 544 -151
rect 823 -145 851 333
rect 540 -169 551 -152
rect 823 -163 829 -145
rect 846 -163 851 -145
rect 517 -188 544 -169
rect 824 -181 851 -163
<< labels >>
flabel metal1 645 265 699 294 0 FreeSans 152 0 0 0 vdd
flabel locali 784 149 813 163 0 FreeSans 104 0 0 0 qbar
flabel locali 551 113 575 128 0 FreeSans 104 0 0 0 q
flabel metal1 646 -43 681 -26 0 FreeSans 120 0 0 0 gnd
flabel locali 545 -168 569 -153 0 FreeSans 120 0 0 0 bl
flabel locali 771 -163 816 -146 0 FreeSans 120 0 0 0 blbar
flabel locali 664 -207 679 -193 0 FreeSans 72 0 0 0 wl
<< end >>
