** sch_path: /home/om/test_first_project/xschem-src/Inverter1.sch
**.subckt Inverter1
Vcc Vcc GND 1.8
vin vin GND pulse(0 1.8 1ns 1ns 1ns 5ns 10ns)
XM1 Vout vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout vin Vcc Vcc sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

 .lib /home/om/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 0.1n  100n
.save all


**** end user architecture code
**.ends
.GLOBAL GND
.end
