magic
tech sky130A
timestamp 1729279079
<< nwell >>
rect 351 381 831 578
<< nmos >>
rect 418 265 433 307
rect 582 265 597 307
rect 722 268 737 323
rect 867 307 909 322
<< pmos >>
rect 418 415 433 457
rect 582 415 597 457
rect 722 402 737 457
<< ndiff >>
rect 680 307 722 323
rect 375 286 418 307
rect 375 269 382 286
rect 399 269 418 286
rect 375 265 418 269
rect 433 303 476 307
rect 433 286 450 303
rect 467 286 476 303
rect 433 265 476 286
rect 539 286 582 307
rect 539 269 547 286
rect 564 269 582 286
rect 539 265 582 269
rect 597 303 640 307
rect 597 286 615 303
rect 632 286 640 303
rect 597 265 640 286
rect 680 290 689 307
rect 706 290 722 307
rect 680 268 722 290
rect 737 307 781 323
rect 867 360 909 364
rect 867 343 878 360
rect 895 343 909 360
rect 867 322 909 343
rect 737 290 754 307
rect 771 290 781 307
rect 737 268 781 290
rect 867 285 909 307
rect 867 268 881 285
rect 898 268 909 285
rect 867 263 909 268
<< pdiff >>
rect 375 442 418 457
rect 375 425 382 442
rect 399 425 418 442
rect 375 415 418 425
rect 433 445 476 457
rect 433 428 449 445
rect 466 428 476 445
rect 433 415 476 428
rect 539 443 582 457
rect 539 426 547 443
rect 564 426 582 443
rect 539 415 582 426
rect 597 443 640 457
rect 597 426 613 443
rect 630 426 640 443
rect 597 415 640 426
rect 680 430 722 457
rect 680 413 688 430
rect 705 413 722 430
rect 680 402 722 413
rect 737 444 781 457
rect 737 430 782 444
rect 737 413 759 430
rect 776 413 782 430
rect 737 402 782 413
<< ndiffc >>
rect 382 269 399 286
rect 450 286 467 303
rect 547 269 564 286
rect 615 286 632 303
rect 689 290 706 307
rect 878 343 895 360
rect 754 290 771 307
rect 881 268 898 285
<< pdiffc >>
rect 382 425 399 442
rect 449 428 466 445
rect 547 426 564 443
rect 613 426 630 443
rect 688 413 705 430
rect 759 413 776 430
<< psubdiff >>
rect 374 166 408 183
rect 425 166 443 183
rect 491 166 515 183
rect 532 166 571 183
rect 830 167 846 184
rect 863 167 910 184
<< nsubdiff >>
rect 375 541 416 558
rect 433 541 448 558
rect 509 541 522 558
rect 539 541 573 558
<< psubdiffcont >>
rect 408 166 425 183
rect 515 166 532 183
rect 846 167 863 184
<< nsubdiffcont >>
rect 416 541 433 558
rect 522 541 539 558
<< poly >>
rect 712 498 747 504
rect 712 481 722 498
rect 739 481 747 498
rect 418 457 433 470
rect 582 457 597 470
rect 712 469 747 481
rect 722 457 737 469
rect 418 371 433 415
rect 582 374 597 415
rect 722 392 737 402
rect 722 377 854 392
rect 388 363 433 371
rect 388 346 396 363
rect 413 346 433 363
rect 388 338 433 346
rect 552 366 597 374
rect 552 349 559 366
rect 576 349 597 366
rect 552 341 597 349
rect 418 307 433 338
rect 582 307 597 341
rect 722 323 737 337
rect 839 322 854 377
rect 839 307 867 322
rect 909 307 922 322
rect 418 252 433 265
rect 582 252 597 265
rect 722 255 737 268
rect 712 247 747 255
rect 712 230 721 247
rect 738 230 747 247
rect 712 220 747 230
<< polycont >>
rect 722 481 739 498
rect 396 346 413 363
rect 559 349 576 366
rect 721 230 738 247
<< locali >>
rect 375 541 383 558
rect 400 541 416 558
rect 433 541 448 558
rect 509 541 522 558
rect 539 541 545 558
rect 562 541 573 558
rect 383 457 400 541
rect 545 457 562 541
rect 712 498 747 504
rect 712 481 722 498
rect 739 481 747 498
rect 712 469 747 481
rect 375 442 410 457
rect 375 425 382 442
rect 399 425 410 442
rect 375 415 410 425
rect 441 445 476 457
rect 441 428 449 445
rect 466 428 476 445
rect 441 415 476 428
rect 539 443 574 457
rect 539 426 547 443
rect 564 426 574 443
rect 539 415 574 426
rect 605 443 640 457
rect 605 426 613 443
rect 630 426 640 443
rect 605 415 640 426
rect 680 430 715 444
rect 459 407 476 415
rect 616 407 633 415
rect 680 413 688 430
rect 705 413 715 430
rect 680 402 715 413
rect 747 430 782 444
rect 747 413 759 430
rect 776 413 782 430
rect 747 402 782 413
rect 388 363 418 371
rect 369 346 396 363
rect 413 346 418 363
rect 388 338 418 346
rect 552 366 582 374
rect 552 349 559 366
rect 576 349 582 366
rect 552 341 582 349
rect 690 364 707 402
rect 459 307 476 313
rect 690 323 707 347
rect 759 364 776 402
rect 759 360 936 364
rect 759 347 878 360
rect 759 323 776 347
rect 867 343 878 347
rect 895 347 936 360
rect 895 343 909 347
rect 867 339 909 343
rect 616 307 633 314
rect 680 307 715 323
rect 441 303 476 307
rect 375 286 410 294
rect 375 269 382 286
rect 399 269 410 286
rect 441 286 450 303
rect 467 286 476 303
rect 605 303 640 307
rect 441 282 476 286
rect 539 286 574 290
rect 375 265 410 269
rect 539 269 547 286
rect 564 269 574 286
rect 605 286 615 303
rect 632 286 640 303
rect 605 282 640 286
rect 680 290 689 307
rect 706 290 715 307
rect 680 281 715 290
rect 746 307 781 323
rect 746 290 754 307
rect 771 290 781 307
rect 746 281 781 290
rect 867 285 909 288
rect 539 265 574 269
rect 867 268 881 285
rect 898 268 909 285
rect 382 183 399 265
rect 547 183 564 265
rect 867 263 909 268
rect 712 247 747 255
rect 712 230 721 247
rect 738 230 747 247
rect 712 220 747 230
rect 875 184 892 263
rect 374 166 382 183
rect 399 166 408 183
rect 425 166 443 183
rect 491 166 515 183
rect 532 166 547 183
rect 564 166 571 183
rect 830 167 846 184
rect 863 167 875 184
rect 892 167 910 184
<< viali >>
rect 383 541 400 558
rect 545 541 562 558
rect 722 481 739 498
rect 459 390 476 407
rect 616 390 633 407
rect 559 349 576 366
rect 690 347 707 364
rect 459 313 476 331
rect 616 314 633 331
rect 721 230 738 247
rect 382 166 399 183
rect 547 166 564 183
rect 875 167 892 184
<< metal1 >>
rect 372 558 573 564
rect 372 541 383 558
rect 400 541 545 558
rect 562 541 573 558
rect 372 535 573 541
rect 712 498 747 520
rect 712 481 722 498
rect 739 481 747 498
rect 712 469 747 481
rect 453 407 482 414
rect 453 390 459 407
rect 476 390 482 407
rect 453 375 482 390
rect 610 407 639 413
rect 610 390 616 407
rect 633 390 639 407
rect 453 366 581 375
rect 453 349 559 366
rect 576 349 581 366
rect 453 341 581 349
rect 610 370 639 390
rect 610 364 714 370
rect 610 347 690 364
rect 707 347 714 364
rect 610 341 714 347
rect 453 331 482 341
rect 453 313 459 331
rect 476 313 482 331
rect 453 307 482 313
rect 610 331 639 341
rect 610 314 616 331
rect 633 314 639 331
rect 610 308 639 314
rect 709 247 766 253
rect 709 230 721 247
rect 738 230 766 247
rect 709 224 766 230
rect 372 184 917 189
rect 372 183 875 184
rect 372 166 382 183
rect 399 166 547 183
rect 564 167 875 183
rect 892 167 917 184
rect 564 166 917 167
rect 372 160 917 166
<< labels >>
flabel locali 369 347 387 362 0 FreeSans 152 0 0 0 in
flabel locali 774 348 808 363 0 FreeSans 152 0 0 0 out
flabel metal1 432 167 475 182 0 FreeSans 152 0 0 0 gnd
flabel metal1 496 351 513 368 0 FreeSans 120 0 0 0 inb
flabel metal1 644 349 666 362 0 FreeSans 120 0 0 0 out1
flabel metal1 459 541 487 557 0 FreeSans 152 0 0 0 vdd
flabel metal1 749 231 766 248 0 FreeSans 120 0 0 0 en
flabel metal1 721 509 737 518 0 FreeSans 120 0 0 0 enb
<< end >>
