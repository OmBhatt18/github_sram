magic
tech sky130A
timestamp 1729278767
<< nwell >>
rect -146 -59 292 -20
rect -146 -198 293 -59
rect -146 -199 246 -198
<< nmos >>
rect -84 -358 -69 -274
rect 54 -357 69 -273
rect 201 -316 216 -274
rect -10 -481 5 -439
<< pmos >>
rect -85 -176 -70 -92
rect 56 -177 71 -93
rect 201 -171 216 -129
<< ndiff >>
rect -126 -330 -84 -274
rect -126 -352 -118 -330
rect -101 -352 -84 -330
rect -126 -358 -84 -352
rect -69 -280 -27 -274
rect -69 -302 -54 -280
rect -37 -302 -27 -280
rect -69 -358 -27 -302
rect 12 -329 54 -273
rect 12 -351 20 -329
rect 37 -351 54 -329
rect 12 -357 54 -351
rect 69 -329 111 -273
rect 155 -289 201 -274
rect 155 -311 163 -289
rect 180 -311 201 -289
rect 155 -316 201 -311
rect 216 -278 255 -274
rect 216 -300 231 -278
rect 248 -300 255 -278
rect 216 -316 255 -300
rect 69 -351 86 -329
rect 103 -351 111 -329
rect 69 -357 111 -351
rect -52 -453 -10 -439
rect -52 -475 -44 -453
rect -27 -475 -10 -453
rect -52 -481 -10 -475
rect 5 -445 48 -439
rect 5 -467 20 -445
rect 37 -467 48 -445
rect 5 -481 48 -467
<< pdiff >>
rect -128 -137 -85 -92
rect -128 -168 -120 -137
rect -102 -168 -85 -137
rect -128 -176 -85 -168
rect -70 -138 -29 -92
rect -70 -169 -55 -138
rect -37 -169 -29 -138
rect -70 -176 -29 -169
rect 13 -138 56 -93
rect 13 -169 20 -138
rect 38 -169 56 -138
rect 13 -177 56 -169
rect 71 -138 112 -93
rect 71 -169 87 -138
rect 105 -169 112 -138
rect 71 -177 112 -169
rect 158 -137 201 -129
rect 158 -161 164 -137
rect 181 -161 201 -137
rect 158 -171 201 -161
rect 216 -137 257 -129
rect 216 -161 233 -137
rect 250 -161 257 -137
rect 216 -171 257 -161
<< ndiffc >>
rect -118 -352 -101 -330
rect -54 -302 -37 -280
rect 20 -351 37 -329
rect 163 -311 180 -289
rect 231 -300 248 -278
rect 86 -351 103 -329
rect -44 -475 -27 -453
rect 20 -467 37 -445
<< pdiffc >>
rect -120 -168 -102 -137
rect -55 -169 -37 -138
rect 20 -169 38 -138
rect 87 -169 105 -138
rect 164 -161 181 -137
rect 233 -161 250 -137
<< psubdiff >>
rect -28 -541 -8 -524
rect 10 -541 129 -524
rect 146 -541 176 -524
<< nsubdiff >>
rect -120 -61 -83 -44
rect -65 -61 41 -44
rect 59 -61 129 -44
rect 147 -61 183 -44
<< psubdiffcont >>
rect -8 -541 10 -524
rect 129 -541 146 -524
<< nsubdiffcont >>
rect -83 -61 -65 -44
rect 41 -61 59 -44
rect 129 -61 147 -44
<< poly >>
rect -85 -92 -70 -79
rect 56 -93 71 -79
rect -85 -205 -70 -176
rect 201 -129 216 -116
rect 56 -205 71 -177
rect -85 -213 71 -205
rect -85 -220 -55 -213
rect -61 -230 -55 -220
rect -37 -220 71 -213
rect 145 -220 176 -210
rect -37 -230 -31 -220
rect -61 -238 -31 -230
rect 145 -237 151 -220
rect 169 -222 176 -220
rect 201 -222 216 -171
rect 169 -237 216 -222
rect 145 -246 176 -237
rect -84 -274 -69 -261
rect 54 -273 69 -260
rect 201 -274 216 -237
rect 201 -329 216 -316
rect -191 -368 -160 -358
rect -84 -368 -69 -358
rect -191 -385 -183 -368
rect -165 -383 -69 -368
rect 54 -382 69 -357
rect 212 -381 243 -371
rect 212 -382 219 -381
rect -165 -385 -160 -383
rect -191 -394 -160 -385
rect 54 -397 219 -382
rect 212 -398 219 -397
rect 236 -398 243 -381
rect 212 -407 243 -398
rect -130 -430 5 -415
rect -130 -451 -115 -430
rect -10 -439 5 -430
rect -138 -461 -107 -451
rect -138 -478 -132 -461
rect -114 -478 -107 -461
rect -138 -487 -107 -478
rect -10 -494 5 -481
<< polycont >>
rect -55 -230 -37 -213
rect 151 -237 169 -220
rect -183 -385 -165 -368
rect 219 -398 236 -381
rect -132 -478 -114 -461
<< locali >>
rect -120 -61 -114 -44
rect -96 -61 -83 -44
rect -65 -61 17 -44
rect 34 -61 41 -44
rect 59 -61 129 -44
rect 147 -61 164 -44
rect -120 -129 -103 -61
rect -128 -137 -95 -129
rect -128 -168 -120 -137
rect -102 -168 -95 -137
rect -128 -176 -95 -168
rect -61 -138 -29 -129
rect 18 -130 35 -61
rect 165 -129 182 -61
rect -61 -169 -55 -138
rect -37 -169 -29 -138
rect -61 -176 -29 -169
rect 13 -138 45 -130
rect 13 -169 20 -138
rect 38 -169 45 -138
rect -55 -205 -38 -176
rect 13 -177 45 -169
rect 80 -138 112 -130
rect 80 -169 87 -138
rect 105 -169 112 -138
rect 80 -177 112 -169
rect 158 -137 190 -129
rect 158 -161 164 -137
rect 181 -161 190 -137
rect 158 -171 190 -161
rect 225 -137 257 -129
rect 225 -161 233 -137
rect 250 -161 257 -137
rect 225 -171 257 -161
rect -61 -213 -31 -205
rect -61 -230 -55 -213
rect -37 -230 -31 -213
rect -61 -238 -31 -230
rect 86 -224 103 -177
rect 145 -220 176 -210
rect 145 -224 151 -220
rect 86 -237 151 -224
rect 169 -237 176 -220
rect -55 -274 -38 -238
rect 86 -241 176 -237
rect -63 -280 -27 -274
rect -63 -302 -54 -280
rect -37 -302 -27 -280
rect -63 -308 -27 -302
rect 86 -323 103 -241
rect 145 -246 176 -241
rect 231 -220 248 -171
rect 231 -237 262 -220
rect 231 -274 248 -237
rect 221 -278 255 -274
rect 155 -289 192 -282
rect 155 -311 163 -289
rect 180 -311 192 -289
rect 221 -300 231 -278
rect 248 -300 255 -278
rect 221 -308 255 -300
rect 155 -316 192 -311
rect -126 -330 -90 -324
rect -126 -352 -118 -330
rect -101 -352 -90 -330
rect -126 -358 -90 -352
rect 12 -329 48 -323
rect 12 -351 20 -329
rect 37 -351 48 -329
rect 12 -357 48 -351
rect 76 -329 111 -323
rect 76 -351 86 -329
rect 103 -351 111 -329
rect 76 -357 111 -351
rect -191 -367 -160 -358
rect -213 -368 -160 -367
rect -213 -384 -183 -368
rect -191 -385 -183 -384
rect -165 -385 -160 -368
rect -191 -394 -160 -385
rect -117 -388 -100 -358
rect 20 -388 37 -357
rect -117 -405 37 -388
rect 20 -439 37 -405
rect 12 -445 48 -439
rect -138 -461 -107 -451
rect -138 -478 -132 -461
rect -114 -478 -107 -461
rect -138 -487 -107 -478
rect -52 -453 -16 -447
rect -52 -475 -44 -453
rect -27 -475 -16 -453
rect 12 -467 20 -445
rect 37 -467 48 -445
rect 12 -473 48 -467
rect -52 -481 -16 -475
rect -130 -504 -113 -487
rect -44 -524 -27 -481
rect 162 -524 179 -316
rect 212 -380 243 -371
rect 212 -381 265 -380
rect 212 -398 219 -381
rect 236 -397 265 -381
rect 236 -398 243 -397
rect 212 -407 243 -398
rect -27 -541 -8 -524
rect 10 -541 129 -524
rect 146 -541 162 -524
rect 158 -545 179 -541
<< viali >>
rect -114 -61 -96 -44
rect 17 -61 34 -44
rect 164 -61 182 -44
rect -44 -541 -27 -524
rect 162 -541 179 -524
<< metal1 >>
rect -120 -44 188 -34
rect -120 -61 -114 -44
rect -96 -61 17 -44
rect 34 -61 164 -44
rect 182 -61 188 -44
rect -120 -70 188 -61
rect 162 -520 179 -515
rect -61 -524 185 -520
rect -61 -541 -44 -524
rect -27 -541 162 -524
rect 179 -541 185 -524
rect -61 -545 185 -541
rect 158 -547 185 -545
<< labels >>
flabel metal1 -58 -60 -10 -45 0 FreeSans 152 0 0 0 vdd
flabel locali 86 -240 122 -225 0 FreeSans 120 0 0 0 dout1
flabel locali 232 -236 260 -221 0 FreeSans 104 0 0 0 dout
flabel locali 244 -396 264 -381 0 FreeSans 120 0 0 0 bl
flabel locali -212 -383 -193 -368 0 FreeSans 96 0 0 0 blbar
flabel locali -129 -503 -114 -488 0 FreeSans 96 0 0 0 ren
flabel locali -54 -262 -39 -244 0 FreeSans 96 0 0 0 2
flabel locali -24 -404 1 -389 0 FreeSans 96 0 0 0 3
flabel metal1 22 -540 75 -525 0 FreeSans 152 0 0 0 gnd
<< end >>
