* SPICE3 file created from replica_bitcell.ext - technology: sky130A
.SUBCKT replica_cell_1rw bl br wl vdd gnd
X0 q vdd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.168 ps=1.64 w=0.42 l=0.15
X1 vdd q vdd vdd sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.64 as=0.4998 ps=4.9 w=0.42 l=0.15
X2 vdd q gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.168 ps=1.64 w=0.42 l=0.15
X3 q vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.62 as=0.168 ps=1.64 w=0.42 l=0.15
X4 q wl bl gnd sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.1722 ps=1.66 w=0.42 l=0.15
X5 vdd wl br gnd sky130_fd_pr__nfet_01v8 ad=0.1596 pd=1.6 as=0.168 ps=1.64 w=0.42 l=0.15
.ENDS
