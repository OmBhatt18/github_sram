magic
tech sky130A
timestamp 1729278616
<< nwell >>
rect -691 98 671 286
rect -691 93 631 98
rect -691 92 72 93
rect -691 91 -63 92
rect -691 86 -64 91
rect -554 85 -411 86
<< nmos >>
rect -628 -29 -613 13
rect -454 -30 -439 12
rect -290 -30 -275 12
rect -145 -30 -130 12
rect -8 -29 7 13
rect 132 -29 147 13
rect 275 -29 290 13
rect 414 -29 429 13
rect 551 -29 566 13
<< pmos >>
rect -628 113 -613 168
rect -456 113 -441 168
rect -290 113 -275 168
rect -145 113 -130 168
rect -10 113 5 168
rect 134 113 149 168
rect 275 113 290 168
rect 414 113 429 168
rect 551 113 568 168
<< ndiff >>
rect -671 0 -628 13
rect -671 -17 -663 0
rect -646 -17 -628 0
rect -671 -29 -628 -17
rect -613 3 -570 13
rect -613 -14 -596 3
rect -579 -14 -570 3
rect -613 -29 -570 -14
rect -498 3 -454 12
rect -498 -14 -490 3
rect -473 -14 -454 3
rect -498 -30 -454 -14
rect -439 2 -394 12
rect -439 -15 -419 2
rect -402 -15 -394 2
rect -439 -30 -394 -15
rect -333 0 -290 12
rect -333 -17 -325 0
rect -308 -17 -290 0
rect -333 -30 -290 -17
rect -275 3 -229 12
rect -275 -14 -258 3
rect -241 -14 -229 3
rect -275 -30 -229 -14
rect -187 1 -145 12
rect -187 -16 -178 1
rect -161 -16 -145 1
rect -187 -30 -145 -16
rect -130 0 -83 12
rect -130 -17 -110 0
rect -93 -17 -83 0
rect -130 -30 -83 -17
rect -52 2 -8 13
rect -52 -15 -44 2
rect -27 -15 -8 2
rect -52 -29 -8 -15
rect 7 2 52 13
rect 7 -15 27 2
rect 44 -15 52 2
rect 7 -29 52 -15
rect 90 3 132 13
rect 90 -14 97 3
rect 114 -14 132 3
rect 90 -29 132 -14
rect 147 1 194 13
rect 147 -16 170 1
rect 187 -16 194 1
rect 147 -29 194 -16
rect 231 0 275 13
rect 231 -17 240 0
rect 257 -17 275 0
rect 231 -29 275 -17
rect 290 3 335 13
rect 290 -14 307 3
rect 324 -14 335 3
rect 290 -29 335 -14
rect 370 0 414 13
rect 370 -17 379 0
rect 396 -17 414 0
rect 370 -29 414 -17
rect 429 3 474 13
rect 429 -14 446 3
rect 463 -14 474 3
rect 429 -29 474 -14
rect 509 3 551 13
rect 509 -14 516 3
rect 533 -14 551 3
rect 509 -29 551 -14
rect 566 2 613 13
rect 566 -15 589 2
rect 606 -15 613 2
rect 566 -29 613 -15
<< pdiff >>
rect -673 144 -628 168
rect -673 124 -665 144
rect -647 124 -628 144
rect -673 113 -628 124
rect -613 144 -569 168
rect -613 124 -593 144
rect -575 124 -569 144
rect -613 113 -569 124
rect -498 151 -456 168
rect -498 121 -491 151
rect -473 121 -456 151
rect -498 113 -456 121
rect -441 151 -394 168
rect -441 121 -420 151
rect -402 121 -394 151
rect -441 113 -394 121
rect -335 151 -290 168
rect -335 121 -328 151
rect -310 121 -290 151
rect -335 113 -290 121
rect -275 151 -231 168
rect -275 121 -258 151
rect -240 121 -231 151
rect -275 113 -231 121
rect -187 152 -145 168
rect -187 122 -179 152
rect -161 122 -145 152
rect -187 113 -145 122
rect -130 151 -83 168
rect -130 121 -109 151
rect -91 121 -83 151
rect -130 113 -83 121
rect -54 151 -10 168
rect -54 121 -47 151
rect -29 121 -10 151
rect -54 113 -10 121
rect 5 159 50 168
rect 5 151 52 159
rect 5 121 26 151
rect 44 121 52 151
rect 5 113 52 121
rect 90 151 134 168
rect 90 121 97 151
rect 115 121 134 151
rect 90 113 134 121
rect 149 151 194 168
rect 149 121 170 151
rect 188 121 194 151
rect 149 113 194 121
rect 230 151 275 168
rect 230 121 238 151
rect 256 121 275 151
rect 230 113 275 121
rect 290 151 334 168
rect 290 121 308 151
rect 326 121 334 151
rect 290 113 334 121
rect 369 151 414 168
rect 369 121 378 151
rect 396 121 414 151
rect 369 113 414 121
rect 429 151 473 168
rect 429 121 448 151
rect 466 121 473 151
rect 429 113 473 121
rect 509 151 551 168
rect 509 121 515 151
rect 533 121 551 151
rect 509 113 551 121
rect 568 151 613 168
rect 568 121 588 151
rect 606 121 613 151
rect 568 113 613 121
<< ndiffc >>
rect -663 -17 -646 0
rect -596 -14 -579 3
rect -490 -14 -473 3
rect -419 -15 -402 2
rect -325 -17 -308 0
rect -258 -14 -241 3
rect -178 -16 -161 1
rect -110 -17 -93 0
rect -44 -15 -27 2
rect 27 -15 44 2
rect 97 -14 114 3
rect 170 -16 187 1
rect 240 -17 257 0
rect 307 -14 324 3
rect 379 -17 396 0
rect 446 -14 463 3
rect 516 -14 533 3
rect 589 -15 606 2
<< pdiffc >>
rect -665 124 -647 144
rect -593 124 -575 144
rect -491 121 -473 151
rect -420 121 -402 151
rect -328 121 -310 151
rect -258 121 -240 151
rect -179 122 -161 152
rect -109 121 -91 151
rect -47 121 -29 151
rect 26 121 44 151
rect 97 121 115 151
rect 170 121 188 151
rect 238 121 256 151
rect 308 121 326 151
rect 378 121 396 151
rect 448 121 466 151
rect 515 121 533 151
rect 588 121 606 151
<< psubdiff >>
rect -674 -107 -640 -90
rect -623 -107 -304 -90
rect -287 -107 -208 -90
rect -191 -107 266 -90
rect 283 -107 343 -90
rect 360 -107 411 -90
<< nsubdiff >>
rect -672 251 -638 268
rect -621 251 -304 268
rect -287 251 -154 268
rect -137 251 264 268
rect 281 251 403 268
rect 420 251 434 268
<< psubdiffcont >>
rect -640 -107 -623 -90
rect -304 -107 -287 -90
rect -208 -107 -191 -90
rect 266 -107 283 -90
rect 343 -107 360 -90
<< nsubdiffcont >>
rect -638 251 -621 268
rect -304 251 -287 268
rect -154 251 -137 268
rect 264 251 281 268
rect 403 251 420 268
<< poly >>
rect -146 215 -115 223
rect -146 198 -139 215
rect -122 198 -115 215
rect -628 180 -441 195
rect -146 187 -115 198
rect -628 168 -613 180
rect -456 168 -441 180
rect -290 168 -275 181
rect -145 168 -130 187
rect -10 168 5 181
rect 134 168 149 181
rect 275 168 290 182
rect 414 168 429 181
rect 551 176 649 191
rect 551 168 568 176
rect -684 52 -649 60
rect -684 35 -676 52
rect -659 50 -649 52
rect -628 50 -613 113
rect -456 100 -441 113
rect -346 76 -311 84
rect -346 59 -338 76
rect -321 74 -311 76
rect -290 74 -275 113
rect -321 59 -275 74
rect -659 35 -613 50
rect -684 29 -649 35
rect -628 13 -613 35
rect -463 49 -428 58
rect -346 53 -311 59
rect -463 32 -455 49
rect -438 32 -428 49
rect -463 25 -428 32
rect -454 12 -439 25
rect -290 12 -275 59
rect -198 74 -167 85
rect -198 57 -192 74
rect -175 73 -167 74
rect -145 73 -130 113
rect -10 84 5 113
rect 134 91 149 113
rect -175 58 -130 73
rect -175 57 -167 58
rect -198 49 -167 57
rect -145 12 -130 58
rect -17 76 13 84
rect -17 59 -11 76
rect 6 59 13 76
rect -17 51 13 59
rect 127 83 157 91
rect 127 66 133 83
rect 150 66 157 83
rect 127 58 157 66
rect 216 76 251 82
rect 216 59 225 76
rect 242 74 251 76
rect 275 74 290 113
rect 242 59 290 74
rect 216 51 251 59
rect -8 13 7 26
rect 132 13 147 26
rect 275 13 290 59
rect 355 76 390 83
rect 355 59 364 76
rect 381 74 390 76
rect 414 74 429 113
rect 551 100 568 113
rect 381 59 429 74
rect 355 52 390 59
rect 414 13 429 59
rect 547 50 577 58
rect 547 33 553 50
rect 570 33 577 50
rect 547 25 577 33
rect 551 13 566 25
rect -628 -64 -613 -29
rect -454 -43 -439 -30
rect -290 -43 -275 -30
rect -145 -43 -130 -30
rect -8 -64 7 -29
rect 132 -64 147 -29
rect 275 -42 290 -29
rect 414 -42 429 -29
rect 551 -42 566 -29
rect 634 -64 649 176
rect -628 -79 649 -64
<< polycont >>
rect -139 198 -122 215
rect -676 35 -659 52
rect -338 59 -321 76
rect -455 32 -438 49
rect -192 57 -175 74
rect -11 59 6 76
rect 133 66 150 83
rect 225 59 242 76
rect 364 59 381 76
rect 553 33 570 50
<< locali >>
rect -672 251 -665 268
rect -648 251 -638 268
rect -621 251 -327 268
rect -310 251 -304 268
rect -287 251 -182 268
rect -165 251 -154 268
rect -137 251 238 268
rect 255 251 264 268
rect 281 251 377 268
rect 394 251 403 268
rect 420 251 434 268
rect -665 155 -648 251
rect -327 159 -310 251
rect -182 159 -165 251
rect -146 215 -115 223
rect -146 198 -139 215
rect -122 198 -115 215
rect -146 187 -115 198
rect 90 159 107 195
rect 238 159 255 251
rect 377 159 394 251
rect -673 144 -639 155
rect -673 124 -665 144
rect -647 124 -639 144
rect -673 113 -639 124
rect -603 144 -569 155
rect -603 124 -593 144
rect -575 124 -569 144
rect -603 113 -569 124
rect -498 151 -467 159
rect -498 121 -491 151
rect -473 121 -467 151
rect -498 113 -467 121
rect -425 151 -394 159
rect -425 121 -420 151
rect -402 121 -394 151
rect -425 113 -394 121
rect -335 151 -301 159
rect -335 121 -328 151
rect -310 121 -301 151
rect -335 113 -301 121
rect -265 151 -231 159
rect -265 121 -258 151
rect -240 121 -231 151
rect -265 113 -231 121
rect -187 152 -153 159
rect -187 122 -179 152
rect -161 122 -153 152
rect -187 113 -153 122
rect -117 151 -83 159
rect -117 121 -109 151
rect -91 121 -83 151
rect -117 113 -83 121
rect -54 151 -23 159
rect -54 121 -47 151
rect -29 121 -23 151
rect -54 113 -23 121
rect 19 151 52 159
rect 19 121 26 151
rect 44 121 52 151
rect 19 113 52 121
rect -739 86 -717 103
rect -700 86 -689 103
rect -684 52 -649 60
rect -708 35 -676 52
rect -659 35 -649 52
rect -684 29 -649 35
rect -597 49 -580 113
rect -498 101 -481 113
rect -546 84 -536 101
rect -519 84 -481 101
rect -597 32 -574 49
rect -557 32 -540 49
rect -597 8 -580 32
rect -498 8 -481 84
rect -411 76 -394 113
rect -346 76 -311 84
rect -411 59 -338 76
rect -321 59 -311 76
rect -463 49 -428 58
rect -463 32 -455 49
rect -438 32 -428 49
rect -463 25 -428 32
rect -411 8 -394 59
rect -346 53 -311 59
rect -259 75 -242 113
rect -198 75 -167 85
rect -259 74 -167 75
rect -259 58 -192 74
rect -259 8 -242 58
rect -198 57 -192 58
rect -175 57 -167 74
rect -198 49 -167 57
rect -111 79 -93 113
rect -52 79 -35 113
rect -111 62 -35 79
rect -111 8 -93 62
rect -52 8 -35 62
rect -17 76 13 84
rect -17 59 -11 76
rect 6 59 13 76
rect -17 51 13 59
rect 35 8 52 113
rect -671 0 -637 8
rect -671 -17 -663 0
rect -646 -17 -637 0
rect -671 -22 -637 -17
rect -603 3 -570 8
rect -603 -14 -596 3
rect -579 -14 -570 3
rect -603 -22 -570 -14
rect -498 3 -465 8
rect -498 -14 -490 3
rect -473 -14 -465 3
rect -498 -22 -465 -14
rect -427 2 -394 8
rect -427 -15 -419 2
rect -402 -15 -394 2
rect -427 -22 -394 -15
rect -333 0 -299 8
rect -333 -17 -325 0
rect -308 -17 -299 0
rect -333 -22 -299 -17
rect -265 3 -232 8
rect -265 -14 -258 3
rect -241 -14 -232 3
rect -265 -22 -232 -14
rect -186 1 -153 8
rect -186 -16 -178 1
rect -161 -16 -153 1
rect -186 -22 -153 -16
rect -119 0 -85 8
rect -119 -17 -110 0
rect -93 -17 -85 0
rect -119 -22 -85 -17
rect -52 2 -19 8
rect -52 -15 -44 2
rect -27 -15 -19 2
rect -52 -22 -19 -15
rect 19 2 52 8
rect 19 -15 27 2
rect 44 -15 52 2
rect 19 -22 52 -15
rect 90 151 121 159
rect 90 121 97 151
rect 115 121 121 151
rect 90 113 121 121
rect 163 151 194 159
rect 163 121 170 151
rect 188 121 194 151
rect 163 113 194 121
rect 230 151 264 159
rect 230 121 238 151
rect 256 121 264 151
rect 230 113 264 121
rect 300 151 334 159
rect 300 121 308 151
rect 326 121 334 151
rect 300 113 334 121
rect 369 151 403 159
rect 369 121 378 151
rect 396 121 403 151
rect 369 113 403 121
rect 439 151 473 159
rect 439 121 448 151
rect 466 121 473 151
rect 439 113 473 121
rect 509 151 540 159
rect 509 121 515 151
rect 533 121 540 151
rect 509 113 540 121
rect 582 151 613 159
rect 582 121 588 151
rect 606 121 613 151
rect 582 113 613 121
rect 90 8 107 113
rect 127 83 157 91
rect 127 66 133 83
rect 150 66 157 83
rect 127 58 157 66
rect 177 76 194 113
rect 216 76 251 82
rect 177 59 225 76
rect 242 59 251 76
rect 177 8 194 59
rect 216 51 251 59
rect 306 76 323 113
rect 355 76 390 83
rect 306 59 364 76
rect 381 59 390 76
rect 306 8 323 59
rect 355 52 390 59
rect 445 77 462 113
rect 509 77 526 113
rect 445 60 526 77
rect 445 8 462 60
rect 509 8 526 60
rect 547 50 577 58
rect 547 33 553 50
rect 570 33 577 50
rect 547 25 577 33
rect 596 8 613 113
rect 90 3 122 8
rect 90 -14 97 3
rect 114 -14 122 3
rect 90 -22 122 -14
rect 162 1 194 8
rect 162 -16 170 1
rect 187 -16 194 1
rect 162 -22 194 -16
rect 232 0 266 8
rect 232 -17 240 0
rect 257 -17 266 0
rect 232 -22 266 -17
rect 300 3 333 8
rect 300 -14 307 3
rect 324 -14 333 3
rect 300 -22 333 -14
rect 371 0 405 8
rect 371 -17 379 0
rect 396 -17 405 0
rect 371 -22 405 -17
rect 439 3 472 8
rect 439 -14 446 3
rect 463 -14 472 3
rect 439 -22 472 -14
rect 509 3 541 8
rect 509 -14 516 3
rect 533 -14 541 3
rect 509 -22 541 -14
rect 581 2 613 8
rect 581 -15 589 2
rect 606 -15 613 2
rect 581 -22 613 -15
rect -665 -90 -648 -22
rect -411 -36 -394 -22
rect -327 -90 -310 -22
rect -179 -90 -162 -22
rect 35 -33 52 -22
rect 35 -52 52 -50
rect 177 -32 194 -22
rect 177 -51 194 -49
rect 238 -90 255 -22
rect 377 -90 394 -22
rect 596 -33 613 -22
rect 596 -54 613 -51
rect -674 -107 -665 -90
rect -648 -107 -640 -90
rect -623 -107 -327 -90
rect -310 -107 -304 -90
rect -287 -107 -208 -90
rect -191 -107 -179 -90
rect -162 -107 238 -90
rect 255 -107 266 -90
rect 283 -107 343 -90
rect 360 -107 377 -90
rect 394 -107 411 -90
<< viali >>
rect -665 251 -648 268
rect -327 251 -310 268
rect -182 251 -165 268
rect 238 251 255 268
rect 377 251 394 268
rect -139 198 -122 215
rect 90 195 107 212
rect -717 86 -700 103
rect -536 84 -519 101
rect -574 32 -557 49
rect -455 32 -438 49
rect -11 59 6 76
rect 133 66 150 83
rect 553 33 570 50
rect -411 -53 -394 -36
rect 35 -50 52 -33
rect 177 -49 194 -32
rect 596 -51 613 -33
rect -665 -107 -648 -90
rect -327 -107 -310 -90
rect -179 -107 -162 -90
rect 238 -107 255 -90
rect 377 -107 394 -90
<< metal1 >>
rect -685 268 434 277
rect -685 251 -665 268
rect -648 251 -327 268
rect -310 251 -182 268
rect -165 251 238 268
rect 255 251 377 268
rect 394 251 434 268
rect -685 240 434 251
rect -685 239 -562 240
rect -151 215 113 223
rect -151 198 -139 215
rect -122 212 113 215
rect -122 198 90 212
rect -151 195 90 198
rect 107 195 113 212
rect -151 189 113 195
rect -723 103 -513 108
rect -723 86 -717 103
rect -700 101 -513 103
rect -700 86 -536 101
rect -723 84 -536 86
rect -519 84 -513 101
rect -723 77 -513 84
rect -20 76 17 84
rect -20 59 -11 76
rect 6 59 17 76
rect 124 83 161 86
rect 124 66 133 83
rect 150 66 161 83
rect 124 59 161 66
rect -580 50 578 59
rect -580 49 553 50
rect -580 32 -574 49
rect -557 32 -455 49
rect -438 33 553 49
rect 570 33 578 50
rect -438 32 578 33
rect -580 25 578 32
rect -419 -33 61 -28
rect -419 -36 35 -33
rect -419 -53 -411 -36
rect -394 -50 35 -36
rect 52 -50 61 -33
rect -394 -53 61 -50
rect -419 -56 61 -53
rect 171 -32 619 -26
rect 171 -49 177 -32
rect 194 -33 619 -32
rect 194 -49 596 -33
rect 171 -51 596 -49
rect 613 -51 619 -33
rect 171 -54 619 -51
rect -679 -90 411 -84
rect -679 -107 -665 -90
rect -648 -107 -327 -90
rect -310 -107 -179 -90
rect -162 -107 238 -90
rect 255 -107 377 -90
rect 394 -107 411 -90
rect -679 -115 411 -107
<< labels >>
flabel locali -597 32 -579 49 0 FreeSans 72 0 0 0 clkbar
flabel locali -234 58 -216 75 0 FreeSans 80 0 0 0 2
flabel locali -85 62 -68 79 0 FreeSans 80 0 0 0 3
flabel locali 177 59 194 76 0 FreeSans 80 0 0 0 4
flabel locali 471 60 490 77 0 FreeSans 80 0 0 0 5
flabel metal1 -541 252 -484 267 0 FreeSans 152 0 0 0 vdd
flabel metal1 -591 -106 -519 -90 0 FreeSans 152 0 0 0 gnd
flabel locali -738 87 -724 102 0 FreeSans 120 0 0 0 din
flabel locali 306 59 336 76 0 FreeSans 120 0 0 0 Q
flabel locali -707 36 -685 51 0 FreeSans 120 0 0 0 clk
flabel locali -394 59 -364 76 0 FreeSans 120 0 0 0 1
<< end >>
