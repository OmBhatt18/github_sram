magic
tech sky130A
timestamp 1729279942
<< nwell >>
rect 699 207 983 349
<< nmos >>
rect 758 40 773 82
rect 907 40 922 82
rect 713 -101 755 -86
rect 859 -101 901 -86
<< pmos >>
rect 758 227 773 269
rect 907 227 922 269
<< ndiff >>
rect 718 70 758 82
rect 718 52 725 70
rect 742 52 758 70
rect 718 40 758 52
rect 773 70 811 82
rect 773 52 788 70
rect 805 52 811 70
rect 773 40 811 52
rect 867 74 907 82
rect 867 51 872 74
rect 889 51 907 74
rect 867 40 907 51
rect 922 75 960 82
rect 922 52 936 75
rect 953 52 960 75
rect 922 40 960 52
rect 713 -54 755 -48
rect 713 -71 723 -54
rect 744 -71 755 -54
rect 713 -86 755 -71
rect 859 -53 901 -48
rect 859 -70 869 -53
rect 890 -70 901 -53
rect 859 -86 901 -70
rect 713 -118 755 -101
rect 713 -135 722 -118
rect 743 -135 755 -118
rect 859 -115 901 -101
rect 713 -142 755 -135
rect 859 -132 868 -115
rect 889 -132 901 -115
rect 859 -141 901 -132
<< pdiff >>
rect 718 262 758 269
rect 718 234 726 262
rect 743 234 758 262
rect 718 227 758 234
rect 773 263 812 269
rect 773 235 787 263
rect 804 235 812 263
rect 773 227 812 235
rect 867 260 907 269
rect 867 235 875 260
rect 892 235 907 260
rect 867 227 907 235
rect 922 261 961 269
rect 922 236 936 261
rect 953 236 961 261
rect 922 227 961 236
<< ndiffc >>
rect 725 52 742 70
rect 788 52 805 70
rect 872 51 889 74
rect 936 52 953 75
rect 723 -71 744 -54
rect 869 -70 890 -53
rect 722 -135 743 -118
rect 868 -132 889 -115
<< pdiffc >>
rect 726 234 743 262
rect 787 235 804 263
rect 875 235 892 260
rect 936 236 953 261
<< psubdiff >>
rect 859 4 884 6
rect 719 -15 761 4
rect 784 -15 823 4
rect 846 -15 907 4
rect 859 -18 884 -15
<< nsubdiff >>
rect 718 300 757 324
rect 781 300 840 324
rect 864 300 909 324
<< psubdiffcont >>
rect 761 -15 784 4
rect 823 -15 846 4
<< nsubdiffcont >>
rect 757 300 781 324
rect 840 300 864 324
<< poly >>
rect 758 269 773 284
rect 907 269 922 284
rect 758 192 773 227
rect 837 194 868 203
rect 837 192 844 194
rect 758 177 844 192
rect 863 177 868 194
rect 758 82 773 177
rect 837 168 868 177
rect 835 134 867 142
rect 907 134 922 227
rect 835 117 842 134
rect 860 119 922 134
rect 860 117 867 119
rect 835 109 867 117
rect 907 82 922 119
rect 758 27 773 40
rect 907 27 922 40
rect 697 -101 713 -86
rect 755 -101 859 -86
rect 901 -101 914 -86
rect 804 -128 819 -101
rect 796 -136 827 -128
rect 796 -153 803 -136
rect 821 -153 827 -136
rect 796 -161 827 -153
<< polycont >>
rect 844 177 863 194
rect 842 117 860 134
rect 803 -153 821 -136
<< locali >>
rect 714 324 909 329
rect 714 323 757 324
rect 714 299 725 323
rect 749 300 757 323
rect 781 300 840 324
rect 864 323 909 324
rect 864 300 871 323
rect 749 299 871 300
rect 895 318 909 323
rect 895 301 953 318
rect 895 299 909 301
rect 714 293 909 299
rect 726 269 743 293
rect 875 269 892 293
rect 936 269 953 301
rect 718 262 751 269
rect 718 234 726 262
rect 743 234 751 262
rect 718 227 751 234
rect 779 263 812 269
rect 779 235 787 263
rect 804 235 812 263
rect 779 227 812 235
rect 867 260 900 269
rect 867 235 875 260
rect 892 235 900 260
rect 867 227 900 235
rect 928 261 961 269
rect 928 236 936 261
rect 953 236 961 261
rect 928 227 961 236
rect 789 159 806 227
rect 837 194 868 203
rect 936 194 953 227
rect 837 177 844 194
rect 863 177 953 194
rect 837 168 868 177
rect 668 142 806 159
rect 668 -56 685 142
rect 789 134 806 142
rect 835 134 867 142
rect 789 117 842 134
rect 860 117 867 134
rect 789 82 806 117
rect 835 109 867 117
rect 936 82 953 177
rect 718 70 749 82
rect 718 52 725 70
rect 742 52 749 70
rect 718 40 749 52
rect 780 70 811 82
rect 780 52 788 70
rect 805 52 811 70
rect 780 40 811 52
rect 867 74 898 82
rect 867 51 872 74
rect 889 51 898 74
rect 867 40 898 51
rect 929 75 960 82
rect 929 52 936 75
rect 953 52 960 75
rect 929 40 960 52
rect 732 12 749 40
rect 873 17 890 40
rect 873 12 907 17
rect 707 7 907 12
rect 707 -17 726 7
rect 751 6 907 7
rect 751 4 864 6
rect 751 -15 761 4
rect 784 -15 823 4
rect 846 -15 864 4
rect 751 -17 864 -15
rect 707 -18 864 -17
rect 889 -18 907 6
rect 707 -22 907 -18
rect 713 -54 755 -48
rect 713 -56 723 -54
rect 668 -71 723 -56
rect 744 -71 755 -54
rect 668 -73 755 -71
rect 713 -78 755 -73
rect 859 -50 901 -48
rect 937 -50 954 40
rect 859 -53 954 -50
rect 859 -70 869 -53
rect 890 -67 954 -53
rect 890 -70 901 -67
rect 859 -75 901 -70
rect 658 -121 683 -112
rect 658 -139 663 -121
rect 680 -122 683 -121
rect 713 -118 755 -112
rect 713 -122 722 -118
rect 680 -135 722 -122
rect 743 -135 755 -118
rect 859 -115 901 -109
rect 680 -139 755 -135
rect 658 -149 683 -139
rect 713 -142 755 -139
rect 796 -136 827 -128
rect 796 -153 803 -136
rect 821 -153 827 -136
rect 859 -132 868 -115
rect 889 -116 901 -115
rect 965 -115 990 -105
rect 965 -116 969 -115
rect 889 -132 969 -116
rect 859 -133 969 -132
rect 986 -133 990 -115
rect 859 -141 901 -133
rect 965 -142 990 -133
rect 796 -161 827 -153
rect 803 -183 821 -161
<< viali >>
rect 725 299 749 323
rect 871 299 895 323
rect 726 -17 751 7
rect 864 -18 889 6
rect 663 -139 680 -121
rect 969 -133 986 -115
<< metal1 >>
rect 657 -121 684 361
rect 708 323 909 336
rect 708 299 725 323
rect 749 299 871 323
rect 895 299 909 323
rect 708 289 909 299
rect 707 7 907 17
rect 707 -17 726 7
rect 751 6 907 7
rect 751 -17 864 6
rect 707 -18 864 -17
rect 889 -18 907 6
rect 707 -25 907 -18
rect 657 -139 663 -121
rect 680 -122 684 -121
rect 963 -115 991 363
rect 680 -139 691 -122
rect 963 -133 969 -115
rect 986 -133 991 -115
rect 657 -158 684 -139
rect 964 -151 991 -133
<< labels >>
flabel locali 804 -177 819 -163 0 FreeSans 72 0 0 0 wl
flabel locali 911 -133 956 -116 0 FreeSans 120 0 0 0 blbar
flabel locali 685 -138 709 -123 0 FreeSans 120 0 0 0 bl
flabel metal1 786 -13 821 4 0 FreeSans 120 0 0 0 gnd
flabel locali 691 143 715 158 0 FreeSans 104 0 0 0 q
flabel metal1 785 295 839 324 0 FreeSans 152 0 0 0 vdd
<< end >>
